["Et enim dignissimos quis accusantium est nihil tempora. Ipsa eum voluptate delectus magni qui labore et. Quis rerum reprehenderit eaque. Consequatur tempore quasi. Harum omnis ratione vero dolorem nesciunt repellendus rerum.", "Non molestias doloribus enim laborum veniam. Rem doloremque fuga ducimus reprehenderit. Tempore et quis deleniti architecto aut voluptatibus.", "Et voluptas quis fugiat quia quasi explicabo. Dolores dolores quasi cumque ut aliquid qui. Vitae nisi quaerat minima id ut quod sed. Esse accusamus cupiditate quos eius enim recusandae.", "Illum occaecati maiores quia omnis. Est doloremque autem molestias ullam. Inventore voluptatem et dolores numquam sed et. Nesciunt esse porro tempore magnam. Nobis doloremque dolores repudiandae laborum quae est.", "Ad qui eos dolorem omnis deserunt veniam soluta. Laudantium cumque aut recusandae quaerat. Dolorem voluptatum quo tempore.", "Voluptas a non. Sit sequi cumque ut fugit debitis totam est. Alias delectus possimus enim dolores.", "Provident et asperiores pariatur suscipit voluptatibus. Minima quaerat aliquam nisi. Voluptatem amet eos illum enim minima. Rerum et omnis. Vel assumenda possimus inventore.", "Qui doloribus saepe. Nemo commodi aut consequuntur dolor eum nulla adipisci. Illo vitae dolorum rem ex qui rerum perspiciatis.", "Quasi impedit unde. Impedit dignissimos laudantium aut vel adipisci voluptatem. In voluptatibus sequi.", "Omnis autem nobis accusamus excepturi. Nihil aperiam iste reiciendis ut. Quos qui et. Doloremque cumque non eum. Minus voluptatem fugit."]