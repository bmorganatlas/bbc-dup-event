["Omnis nulla at ipsam. Quis iure autem est molestias qui. Tempora qui ad laboriosam culpa occaecati non distinctio.", "Omnis modi dolorum voluptatem optio. Et eos magnam placeat quae accusantium sint accusamus. Error et tenetur ut debitis fugit. Atque ab quis aut maxime commodi. Et numquam corrupti dignissimos dolores vitae exercitationem et.", "Laudantium commodi adipisci voluptatem tenetur vel. Veritatis laborum sapiente eligendi at voluptatum. At magnam vel expedita odit. Reprehenderit fugiat ut.", "Sequi qui aut eveniet. Aut fugit ea. Eveniet quia reprehenderit assumenda vero quasi aliquid. Quas doloremque at voluptatibus et commodi est. Odio nisi est vero dicta molestias neque tempora."]