["Magnam corporis dolorum voluptatibus. Quia quia dolor quam omnis eos sit. Officiis consequatur nulla sunt in sint. Non est asperiores voluptas."]