["Quasi ducimus dicta neque fuga quia. Dolorem ipsam occaecati. Quaerat ut natus blanditiis voluptatem placeat quod sit."]