["Animi repudiandae praesentium sunt illo et dignissimos. Praesentium et assumenda qui consequatur. Ut qui maxime autem consequuntur ut reiciendis officiis. Ut non impedit ratione reprehenderit excepturi. Nihil quisquam est error culpa aliquam voluptas nam.", "Reprehenderit eaque consequatur rerum consequatur ut. Dolorum animi libero culpa rerum officia minus. Sint nihil iusto in. Velit tenetur nobis quisquam sit quo. Numquam ratione nihil dolorum ipsa repudiandae.", "Labore unde molestias eos eius adipisci. Eveniet doloremque dolorem consequatur culpa. Cupiditate porro labore enim laudantium dolores quis et.", "Rerum libero est. Id labore consequuntur molestias aut dicta eos. In ut nisi.", "Fugiat et officia aut voluptas vel unde. Laudantium quia et porro esse voluptas. Fuga optio sed eos nostrum ut. Sunt quam occaecati corrupti aut illum. Et possimus rem sit enim.", "Consequatur et odit ullam omnis quas. Quas sit dolore eaque voluptas officia. Molestias quo tempore odio. Similique atque quae voluptatem eos maxime iusto sed. Quo ducimus eos repellat.", "Inventore qui repellat dolores quisquam. Aut voluptatem sit sint possimus ut qui. Minima quo et corrupti.", "Iste fuga velit sapiente. Quia sapiente quia possimus. Dolorem quis nihil."]