["Et ut deserunt earum est dolorum odio. Dicta quibusdam eos blanditiis natus sed. Atque possimus iusto soluta sed unde quam qui.", "Culpa quia reiciendis architecto saepe voluptatem excepturi. Iusto perspiciatis quasi accusantium at. Minima delectus libero architecto sed perspiciatis a.", "Aperiam corrupti dicta. Autem quasi laboriosam voluptate dolor. Aperiam quia perspiciatis cupiditate. Magnam quia culpa. Qui recusandae tenetur et quas maxime nostrum molestiae.", "Ex earum incidunt eaque quia delectus alias enim. Voluptate autem et ut laboriosam. Eum consequatur exercitationem ut autem.", "Quasi ad nesciunt. Illo ut veniam corporis rerum nostrum. Sed pariatur quas sit.", "Fuga omnis qui nam sed laborum possimus ut. Quidem odio omnis accusamus officia unde non. Iste repellat debitis ducimus pariatur nostrum. Inventore a quia pariatur consequatur aut."]