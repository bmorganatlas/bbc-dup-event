["Ex veniam omnis. Ut voluptas occaecati officia. Velit libero dolores reiciendis dolores sint. Tempore quaerat iusto. Dolores vel et.", "Sapiente tempora labore excepturi amet magnam. Aliquam nulla eius provident laborum et. Accusamus non a suscipit dolorem. Perferendis officiis repudiandae voluptatum.", "Deserunt recusandae aut minus delectus omnis. Dolorem sunt ut neque. Ipsam enim voluptatem porro itaque voluptatem.", "Perferendis repellat distinctio voluptas molestias voluptatem quibusdam. Placeat maiores id quae tempore occaecati repudiandae. Ea facere vel non. Et culpa aperiam incidunt officia sint."]