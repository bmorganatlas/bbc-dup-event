["Magni eum quia. Quis quibusdam dolorum aperiam eaque non maiores. Sint eligendi velit maiores.", "Minima eos quia. In earum cum cupiditate molestiae sint aut enim. Ea ipsa omnis itaque sint incidunt perferendis. Quis aliquam nostrum minus asperiores et. Inventore nesciunt veritatis omnis et reiciendis et vel.", "Est est sapiente ducimus esse laborum sunt voluptatum. Qui quas illum et perferendis aut laborum. Voluptate qui dolor soluta error necessitatibus qui.", "Sit sint enim. Et ut rerum assumenda. Omnis repellendus eos assumenda nihil et quis ut. Voluptatem sit velit quo et eum quibusdam nobis.", "Omnis maiores necessitatibus illo. Tempore exercitationem numquam. Consequatur unde dolor aut quos. Autem ipsum tempore non minus. Et veniam velit ea nobis.", "Deserunt eius qui aliquid aut id. Enim et sequi qui rerum nam repellendus. Repellendus laboriosam modi cum. Expedita culpa est officiis.", "Voluptates sit unde tempora aut voluptatem. Fugit cumque saepe ratione sit sapiente est quia. Beatae odit ducimus ea ipsum modi omnis.", "Explicabo eveniet et. Sed quia perferendis fugit consectetur. Fugiat et eius vitae repellendus dolores consequatur maiores. Minus neque nesciunt ipsa a. Voluptatem officiis beatae.", "Incidunt eum impedit. Alias eum nam velit enim. Ad doloribus quae ut. Voluptatem sunt quia natus corrupti. Quidem eligendi eos ea repellat debitis corrupti.", "Consequatur sunt ut dolorum beatae dolorem fugit ab. Tenetur distinctio voluptatum expedita nam quam et. Velit unde ipsam blanditiis laboriosam dolorum. Id atque non et ipsam. Nisi sed a impedit."]