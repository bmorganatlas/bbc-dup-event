["Similique quod consequuntur praesentium unde. Sunt et voluptas voluptas eos. Corrupti illo et commodi.", "In dolorum consequatur. Non qui repellat molestiae alias facere qui quia. Quae soluta reprehenderit corrupti.", "Quia officiis magnam quia molestiae. Ut facilis neque. Dolore quo illum. Iste quas magni delectus doloribus minima. Et eum quo ut fuga veritatis animi possimus.", "Molestiae itaque dolorem nulla praesentium veritatis sit sint. Non odit reprehenderit quia. Adipisci debitis nihil perspiciatis et fugit aut nemo. Accusamus aut ex ducimus sed blanditiis tempore.", "Porro ipsum ullam magnam quo rem. Eligendi molestias laborum et quisquam alias. Velit aut magnam est repellat quibusdam tenetur autem. Qui quo aut consequuntur. Ab sed alias sequi quidem quae nisi.", "Placeat velit ratione et sed aspernatur accusantium. Veritatis consequatur commodi repellat nemo eos ea. Illo eius et dolor. Repellat similique repudiandae vero.", "Sunt id rerum doloribus. Minus qui fugit adipisci molestiae dolores assumenda aut. Quas similique omnis et sed accusantium rerum nostrum.", "Occaecati qui laborum. Et voluptatum beatae velit. Pariatur ut quia quod. Ea in voluptate. Est et maiores est illo ipsa.", "Sapiente voluptate fugit consequatur molestias. Ullam rerum recusandae mollitia ut adipisci. Facilis consectetur illum cumque est blanditiis. Libero eveniet distinctio velit reprehenderit.", "Facere recusandae reiciendis dolore est sed. Aliquid quidem quia veritatis itaque fuga qui sed. Architecto fuga error dignissimos. Itaque aliquam tempora quasi magni quaerat voluptatem."]