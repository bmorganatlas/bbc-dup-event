["Omnis repudiandae quidem et. Voluptatem et voluptate sequi a dolor id aut. Sunt quis aut ipsa reiciendis rerum autem debitis. Quae ut ea nihil omnis enim. Veritatis ex tenetur architecto.", "Voluptatum repudiandae illo alias pariatur. Est quo porro pariatur aut non. Non error dicta repellendus."]