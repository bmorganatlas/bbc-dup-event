["Aut molestiae rem. Totam et possimus. Omnis doloribus quisquam illum veniam.", "Distinctio doloremque non quaerat eius. Dolorem asperiores fugit nihil. Velit incidunt qui quaerat eius atque. Dolor eos et est occaecati quia doloremque quo. Error placeat eos rerum et nulla in molestiae.", "Ea aliquam animi. Iure porro omnis. Dignissimos illum quis aut voluptatem debitis ratione corporis.", "Et nihil doloribus. Quam porro cumque. Est sequi sint qui dolores. Iure voluptas consequatur corrupti aut asperiores ea. Aut officia ex eos iste qui enim.", "Repellendus et ut sit reprehenderit id. Eos libero consequuntur nihil. Iure et ex aut atque et.", "Expedita odit sit. Explicabo possimus sapiente. Ducimus optio aut minus possimus rerum explicabo. Officia ut reprehenderit.", "Voluptatem consequatur quaerat tempora asperiores. Enim ullam sint eveniet vero. Et eveniet placeat illum labore error dolorem. Culpa hic ipsa iste aperiam. Eos quia assumenda harum odit earum qui.", "Ea dolores deleniti. Tempora maiores officia. Alias atque numquam ea veniam praesentium id. Culpa in alias.", "Quam quo impedit aut voluptatem voluptatem nulla. Et qui fuga amet ea rerum. Rerum assumenda labore quas delectus excepturi.", "Delectus beatae eos. Consequuntur distinctio enim. Voluptatem voluptatibus porro reprehenderit nostrum ratione et. Consequatur officiis nostrum officia. Praesentium quia veniam consequatur optio ut."]