["Ut sed nihil. Suscipit exercitationem quis sint. Ipsam sit qui.", "Maxime enim culpa praesentium dolorem ad. Deserunt doloremque pariatur. Qui laborum ut sit. Modi tempore molestiae. Est cumque ea voluptas facilis magnam et laboriosam.", "Dignissimos occaecati mollitia iusto provident et eius ut. Ab atque quis excepturi minima quae. Deleniti voluptates ipsam accusamus vel.", "Beatae assumenda voluptatem harum fugiat asperiores optio. Et numquam nulla tenetur cum quibusdam consequatur aut. Id nostrum aut totam illo velit voluptatem ut. Nesciunt fugit minus praesentium pariatur eveniet. Non sequi sint tempore quis laudantium.", "Fugiat qui et repudiandae iure facilis veritatis quas. Quis incidunt voluptate. Quisquam assumenda maiores excepturi non eaque."]