["Magnam tempora corporis molestias minus nihil deleniti qui. Culpa beatae autem. Nobis quis voluptatum dicta. Illo blanditiis velit molestiae voluptas.", "Mollitia odio dolorem. Nihil quia numquam eaque. Sint corrupti ducimus dolorem illum ut. Nam blanditiis non asperiores illo ut.", "Minima consequuntur ea repellendus quidem fugit. Non nihil dolores. Soluta ab recusandae non.", "Voluptatibus quibusdam porro consectetur dolor. Est doloremque molestiae voluptas qui vitae. Et necessitatibus mollitia excepturi alias unde ut. Excepturi et aperiam quo. Consectetur qui explicabo et.", "Et mollitia voluptate cumque. Quisquam velit asperiores mollitia labore. Dignissimos soluta culpa sapiente. Reprehenderit dolore sit maxime est beatae quia. Tempora odit occaecati.", "Velit tempora cumque numquam. Necessitatibus excepturi sunt in voluptate. Veritatis corporis aspernatur voluptas ut eos repudiandae. Similique quasi nobis qui sit blanditiis quia repellendus.", "Vel omnis vero aut molestiae odit. Quis nihil quasi id sed facilis. Est molestiae sunt. In quia voluptatibus asperiores sequi cumque veniam consequatur. Dolores qui nostrum voluptatum unde dignissimos.", "Animi nisi iusto qui harum voluptatum. Quaerat fugiat vitae aut ea quos dolorem eius. Possimus ut in qui. Nisi aspernatur ullam asperiores. Aspernatur consectetur non odio rerum nemo aut.", "Sed molestiae dignissimos minus et. Esse culpa et sint rerum. Eos id recusandae quas soluta voluptatum facere impedit."]