["Id explicabo eveniet non sed. Consequatur quod dolorem id nihil. Dolores molestiae vero voluptas debitis voluptatem. Architecto id aut aspernatur.", "Qui omnis recusandae non labore repudiandae asperiores et. Rerum pariatur deserunt perferendis et iure. Officiis et optio."]