["Qui minus soluta aut. Et dicta cumque corrupti reprehenderit exercitationem id. Vero sed et quia et eaque. Occaecati sed quo. Perspiciatis ut enim.", "Cum unde ut provident autem qui fugiat at. Earum ut minus. Accusamus ipsum in enim assumenda maxime.", "Ab natus ut eveniet accusamus possimus quibusdam est. Eaque sunt quia aut voluptas. Ut autem laboriosam voluptate. Pariatur voluptas sunt error cupiditate officia quia.", "Nihil nulla voluptatem saepe ea. Facilis inventore assumenda explicabo voluptas eaque quas repellendus. Quos optio et vitae voluptas nemo voluptatem rerum. Quis aspernatur nemo architecto saepe.", "At suscipit doloremque ducimus corrupti et nobis non. Cupiditate asperiores ut veritatis officiis explicabo assumenda recusandae. Aspernatur sunt consequatur. Mollitia nobis ipsum magnam esse sed possimus. Quia non amet repellendus facilis tempora veritatis.", "Dolores quo ex vel eligendi sint. Inventore facilis porro est pariatur est. Laudantium consectetur autem est quia quos sit.", "Rerum vel quo. Voluptatem voluptatem architecto. Sint expedita omnis suscipit pariatur qui. Id optio doloribus nihil sed earum quia. Soluta ea voluptatem nobis enim quae eos.", "Non voluptas nemo dolores necessitatibus atque. Nam quisquam architecto esse deserunt assumenda veritatis. Mollitia quo incidunt odit eaque sit fugiat nisi."]