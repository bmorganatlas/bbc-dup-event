["Dicta placeat consequatur sed rerum blanditiis sunt minus. Sunt libero quis sint reprehenderit quam maiores. Modi aut dolorum aut et sunt.", "Rem aut ipsam enim non incidunt eos. Quasi repellat quisquam vero. Facere aperiam voluptatem repellendus repudiandae ut.", "Culpa quidem officia. Dicta commodi voluptatem. Distinctio quibusdam odit aut temporibus in. Eius sed ipsum ab necessitatibus ea est velit.", "Dolorum dolores qui est. Dolorum inventore consequatur ut. Eos facere vel voluptas et. Explicabo sequi voluptate mollitia."]