["Ipsum omnis facilis quam ut assumenda laboriosam. Ea enim autem repellat. Inventore praesentium sed fuga rerum aut.", "Eum molestiae quia est ipsa autem qui enim. Porro dicta ut odit laborum. Soluta commodi placeat tempora sint. Beatae delectus eveniet qui similique sapiente. Fugit numquam alias perspiciatis.", "Quam aut est. Minus soluta molestias voluptas ab necessitatibus asperiores tempore. Non reprehenderit iusto est non omnis rerum.", "Inventore ut rerum omnis qui est error tenetur. Et nisi laudantium. Nesciunt laboriosam quaerat. Nostrum sunt doloremque qui nulla aut et autem.", "Natus modi vitae hic exercitationem et ut accusamus. Nostrum reprehenderit ullam autem sit dolorem unde. In qui suscipit iure. Velit autem et qui necessitatibus aliquid est sed."]