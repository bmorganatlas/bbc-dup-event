["Ipsa alias odio. Cupiditate vitae quod est qui tenetur et nulla. Est optio fugiat debitis et impedit distinctio. Mollitia quos facere.", "Voluptatem quia dolor nemo qui. Aspernatur laudantium mollitia dolorum. Assumenda rem dolores ratione. Quibusdam unde consequatur. Rerum perspiciatis omnis.", "Sunt voluptas blanditiis qui vitae eligendi est. Velit aliquid sed sequi blanditiis ea exercitationem et. Enim placeat aut unde sunt hic rerum excepturi. Ullam molestiae quo aut illo facilis. Sed odio quasi non atque porro.", "Non fuga et. Aut ad autem eligendi. Fugit explicabo quidem minima.", "Est aperiam reprehenderit. Qui qui in ea sint. Accusantium et aut.", "Aspernatur repudiandae corporis. Laboriosam vel placeat cumque rerum quo et. Nulla culpa esse aspernatur explicabo et. Labore perspiciatis tempora eius autem fugiat vel. Et enim culpa voluptas ullam aliquam iste aut.", "Et quae sequi quis sapiente aut. Sunt ut iure. Vitae ipsa molestiae sit sed deserunt ut.", "A mollitia atque quidem. Ullam aliquid eum ab. Quaerat dignissimos nobis architecto consequatur.", "Possimus sit voluptatum. Nulla officia et corrupti non. Odit reprehenderit sit dolor reiciendis autem in.", "Deserunt asperiores omnis. Repellat corrupti consequuntur voluptas. Est nobis ipsum. Qui sunt quo hic expedita."]