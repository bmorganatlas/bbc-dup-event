["Aspernatur consequuntur repudiandae dolores. Molestias aspernatur doloremque assumenda et. Voluptas hic est dolorum quidem consequatur incidunt dolorem.", "Occaecati omnis temporibus et praesentium nemo ullam. Vitae odit et iste ea et. In et voluptatem expedita possimus omnis. Possimus ut nobis facilis.", "Dolor reprehenderit autem qui et mollitia asperiores officiis. Error in nemo voluptas consequatur. Consequatur exercitationem adipisci iusto. Repudiandae non reiciendis ex eligendi. Magni enim eveniet quisquam facere quae.", "Quasi debitis totam. Adipisci enim amet. Sed temporibus distinctio.", "Libero veritatis dolore sit sint omnis consequatur. Deserunt asperiores soluta amet tempora est. Veritatis delectus autem reiciendis voluptate et id. Qui voluptates ut ut. Labore ut omnis.", "Distinctio aut tempora nisi adipisci earum ut quisquam. Aut facere totam voluptas consequatur dolore. Qui magni sint. Velit minus aliquid placeat earum fuga rerum."]