["Ut et cumque. Tenetur cum voluptatem qui. Praesentium dicta commodi veniam nobis modi ad. Ipsam consequuntur enim quasi eius suscipit. Ut voluptatum error.", "Molestias nesciunt fugit enim. Quod earum aperiam molestiae tenetur. A corporis veritatis dolorum quo dignissimos. Molestias fuga rerum expedita. Eaque quam quis.", "Praesentium et nam. Qui hic ut vel ut in voluptatum ipsa. Omnis voluptatem et adipisci natus amet quia molestiae.", "Quae earum ea voluptates eligendi sint sed. Odio tenetur velit sed dignissimos ut. Laborum aut nihil. Itaque numquam eius natus maiores et ut. Nostrum vitae optio.", "Ratione voluptate sint. Iusto iure assumenda vero. Voluptatem velit quia corrupti commodi nulla. Similique dolorem quia.", "Enim omnis maiores ut. Ipsum cum dolor cumque. Minima asperiores quia officia eligendi. Est suscipit laboriosam."]