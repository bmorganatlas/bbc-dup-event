["Ratione aut qui. Libero rerum minima in. Officia vel molestiae. Veniam mollitia sint recusandae.", "Eum dolores sequi praesentium ipsum aliquam voluptates. Sed provident dolor necessitatibus distinctio occaecati amet molestiae. Id recusandae fuga.", "Quia perferendis dignissimos. Est eveniet in fugiat reprehenderit sed. Voluptates eum possimus vel sequi accusantium incidunt enim.", "Et pariatur eaque eum earum et quibusdam dolorem. Cum et ducimus minima corporis non pariatur. At fuga eligendi animi blanditiis doloremque est. Excepturi odit aut explicabo sed in ut. Nobis dolorem et.", "Tempore quod sit et voluptatem eveniet. Consectetur necessitatibus ex facilis aut nobis corrupti. Nam ducimus et.", "Aut laudantium consequatur distinctio optio cumque magni. Explicabo accusantium rerum. Dicta id consequatur fugit dolore delectus.", "Ipsam voluptatibus in. Dicta et quis molestiae. Nostrum inventore ad sequi. Qui mollitia quasi ut est libero. Eligendi placeat culpa odio voluptates.", "Et ullam autem eum hic. Provident sunt tenetur vero. Aut voluptatem aperiam.", "Voluptate aut et porro maxime molestiae. Incidunt fugit quod ratione. Quod eveniet sequi dolorum. Sit et ab. Occaecati harum eligendi esse non ut.", "Mollitia qui eveniet et nihil eum quas. Quos est aliquam dolor. Ipsa iusto suscipit voluptates debitis. Pariatur quae earum ad. Dolore autem dolorem neque."]