["Dolor voluptate eaque quasi est aliquid quia. Qui qui quo tenetur. Est eum nesciunt neque cumque occaecati. Natus id nihil molestias.", "Quisquam voluptatem possimus qui sed impedit ut aut. Ut eum et expedita sint maiores vel. Sed nemo ipsam esse.", "Voluptatum tempore ab aut ut. Nulla non corporis sequi. Eos a corrupti sit ab totam maiores voluptatem. Tempora maiores incidunt tempore dicta."]