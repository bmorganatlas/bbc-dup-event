["Numquam eaque eum id consequuntur eligendi hic autem. Blanditiis laudantium fugiat beatae nihil dicta. Placeat officiis nesciunt illum magnam. Similique non adipisci eveniet sed sed. Error et iste sint quibusdam dolores.", "Eos enim vitae. Commodi atque tenetur. Ut et nostrum nemo repudiandae. Laborum reprehenderit quia possimus."]