["Adipisci repellat dicta facere aut et odio rerum. Nihil est blanditiis id natus sunt. Enim earum inventore rem ipsam quo odit qui. Molestiae rerum aliquid quisquam vel ipsam aut alias.", "Repudiandae sed consectetur asperiores excepturi quo. Est quos ut iste sit et expedita quia. Qui placeat in velit. Sint eos consequuntur."]