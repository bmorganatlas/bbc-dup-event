["Deleniti nam perferendis ipsam necessitatibus id velit distinctio. Corrupti dolores distinctio. Libero quas ratione doloremque officiis.", "Sunt minima alias et excepturi dolorem. Consequatur amet ex non autem temporibus omnis. Sint sunt optio aut quia. Est nihil at amet quasi. Fugit illum blanditiis quaerat odio quae.", "Molestiae molestias beatae qui quos voluptatibus pariatur non. Et modi est repudiandae. Odit aperiam doloremque corporis. Illum odio cumque ab voluptatem nulla ipsum tempora. Cum ut ut et unde recusandae aut.", "Sunt est totam cumque dolores rerum libero. Sed quis iusto eum et veniam. Et rerum nemo quos voluptas enim qui sequi. Laboriosam animi cupiditate magnam consequatur. Voluptate omnis autem.", "Voluptas deserunt ipsa. Aut alias natus error qui sit quam. Sunt in eos aliquam. Aperiam optio vel sed.", "Minus nisi tempore porro sit sint est cum. Porro aliquam optio vitae non amet sint nesciunt. Soluta minima non."]