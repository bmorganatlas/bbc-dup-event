["Qui enim cumque eius totam optio quia delectus. Nemo excepturi aspernatur. Accusamus soluta fugit consequatur voluptatum minima. Cumque quaerat ducimus sapiente. Suscipit dolorem occaecati ab.", "Nihil placeat perferendis minus quos quas quo vel. Officia minima ab commodi sed quia. Qui quae voluptas assumenda. Blanditiis est velit sint et. Quis velit qui atque harum.", "Qui praesentium aliquam voluptatem occaecati debitis. Fugit reprehenderit iure eum qui. Est velit vel sunt. Vel quo quis quisquam alias sint excepturi.", "Vel modi nulla ut doloribus eveniet rerum veniam. Architecto eligendi occaecati et voluptatem at. Quia quam soluta rerum ut. Qui harum quae aspernatur vel quasi. Dolor est illum.", "Provident minima officiis. Doloribus modi perspiciatis dolores similique repellendus. Consequatur ut doloremque qui omnis possimus minus. Neque repellendus illum quibusdam ut.", "Ut cupiditate debitis eum quidem corporis et. Dolor culpa cumque aliquid blanditiis voluptatem quasi. Sint consequatur voluptatem in ut. Numquam officiis quia veniam esse dicta ut exercitationem. In necessitatibus eum neque."]