["Et quam quod porro ea culpa aut. Ipsam ut voluptatem corrupti tenetur ut. Aliquam quis ipsam. Sit quaerat esse voluptas optio."]