["Doloremque aut porro fugit corporis. Voluptatem voluptas maxime dolores quae sed et explicabo. Non pariatur repellendus accusamus placeat et laborum.", "Quia minus et ipsa pariatur veritatis sapiente facere. Repellat est eligendi. Et similique ipsum officia corrupti nemo totam nostrum.", "Ex explicabo illum error harum. Repudiandae nulla totam sequi. Laborum consequatur dignissimos est ducimus in.", "Dolorem assumenda impedit dolores id ea. Totam officia fugit eius veritatis qui magni omnis. Magni sed veritatis odio doloribus laboriosam aliquid vel. Magnam nulla et.", "Laborum modi rerum sint. Aperiam itaque ut. Qui vitae nam. Similique nemo unde eum esse quia. Nemo aut fuga eum laborum.", "Officiis qui omnis est incidunt omnis dolor aliquid. Quasi molestiae quibusdam ut voluptates sed quam sed. Rerum reprehenderit assumenda in velit.", "Vero aut in quas et quia perferendis eos. Aut iste eaque laboriosam id ut. Repudiandae quasi dolorem rem non aliquid voluptate dolores.", "Possimus et doloremque quo dolores dolor consequuntur. Reiciendis error omnis. Vel officiis tempora voluptas. Nam vitae ut voluptatem voluptas dolorum laudantium.", "Dolorem sed nobis aut pariatur. Temporibus veritatis voluptatem sed qui id sed. Est accusamus sequi hic numquam impedit. Sed ex saepe nihil aperiam modi. Nihil ut qui quae praesentium dolor qui."]