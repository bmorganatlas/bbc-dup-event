["Quis error ut. Enim sed accusantium non qui ipsum vel. Quos natus aut nihil et laborum repellendus.", "Eaque ab quisquam qui sint asperiores iusto fugit. Enim assumenda officia qui natus debitis iure minima. Et consequuntur magni officiis enim voluptas magnam nesciunt.", "Quidem et ut. Eum veniam unde illum ut. Alias expedita et aut aut consectetur maxime eos.", "Dolorem doloremque aut error quam saepe. Inventore ad et corrupti. In quod atque.", "Quidem perferendis omnis dolorem magnam rem aperiam. Officiis accusamus dolorem sint. Impedit provident explicabo sed. Optio vel et voluptatem dignissimos deleniti. Beatae ipsum repellat nulla incidunt.", "Voluptates dolores odit. Nihil ut reprehenderit est eum quam ipsa. Officia molestiae dolorem. Amet qui nihil et. In eligendi reprehenderit deserunt ut unde sint repellendus.", "Id et aut. Nisi quos corporis. Eum libero incidunt dolorem. Nobis nisi dolorem voluptates repellat et.", "Ullam occaecati corrupti provident vitae. Recusandae veritatis aut vitae dolorem. Rerum modi nulla officiis itaque. Quos iusto et.", "Dicta impedit excepturi. Dolore ullam asperiores quo qui omnis. Sed omnis explicabo ea reprehenderit quidem quibusdam. Culpa illo modi. Architecto rerum harum porro quia expedita repudiandae omnis.", "Aut ut excepturi. Facilis ad sint quod id nemo dolore quidem. Harum ab minima. Omnis minima quidem quam vel maxime ipsa iste. Iste quidem velit."]