["Ab perspiciatis consectetur quisquam quo non. Iusto rerum delectus vero laudantium. Animi aperiam commodi. Illo in voluptatem excepturi accusamus modi. Aut reprehenderit dicta ipsam natus.", "Provident et maxime. Cum enim eos. Maxime debitis recusandae voluptate aliquid.", "Numquam itaque similique saepe. Molestiae quia ut. Adipisci quisquam quia. Quasi et rem deserunt.", "Quasi autem voluptate molestiae. Inventore culpa dolor asperiores quo animi. Ut in odio. Veritatis sequi quia fugit dolores deleniti.", "Quibusdam commodi in. Voluptatem magnam qui autem neque repellendus ipsam. Odio et nam rem est. Magnam molestiae maxime voluptate id earum omnis. Eum dolore maiores sit qui quo dolores eveniet.", "Vel dolor eveniet. Amet eos et. Consequuntur exercitationem dolorem aliquam voluptatibus aspernatur."]