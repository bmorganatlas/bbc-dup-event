["Nihil quia et excepturi. Et officiis ratione tempora non. Voluptatem molestiae voluptatibus quia et. Et optio et sapiente porro animi. Architecto in fugiat ipsum et.", "Sit qui quod dolores temporibus. Aut inventore ex. Libero sunt et consectetur quia. Quae consequatur nobis nostrum voluptatem voluptatum laborum sit. Dolore voluptas incidunt ratione iusto.", "Qui sapiente ipsam autem. Minima illo molestiae harum explicabo. Velit est aperiam. Aut accusamus et. Deleniti corporis aut.", "Deserunt qui illum. Vitae iusto magni necessitatibus quod. Dolor esse dolores.", "Error aut dolorum alias enim nisi tenetur omnis. Quis est rerum autem necessitatibus unde dolorem corporis. Sint pariatur aut ipsa quia adipisci. Itaque et ipsam voluptate odit. Voluptatem natus repellendus et error et.", "Eum maxime assumenda. Beatae et unde asperiores deleniti aut odio. Laborum illum omnis sunt. Voluptas accusantium id.", "Dolores ipsum eaque porro. Harum eos aut. Rerum pariatur odio amet omnis ut impedit.", "Reprehenderit molestiae voluptas. Aut consequatur dolorem. Dolore et perspiciatis et molestias consequatur inventore et."]