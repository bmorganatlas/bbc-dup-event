["Quaerat repellendus alias necessitatibus in. Modi repellendus qui aliquid commodi eius. Rerum incidunt pariatur reiciendis quis. Maiores omnis repellat soluta explicabo consequatur quisquam saepe.", "Beatae molestiae eveniet dignissimos voluptates. Non velit aut. Dignissimos reprehenderit cumque. Unde earum a inventore aperiam. Et deleniti suscipit ut.", "Dolorem nulla qui sunt dolore soluta inventore quis. Ad consequatur aut non quasi velit fugiat. Eaque rem debitis qui sed iusto itaque. Eos et sed.", "At vero voluptatibus. Dolorem similique corrupti cum. Aut qui quis vel quia adipisci.", "Quo ea est. Expedita voluptatem ea ab voluptatem occaecati et. Possimus tempore molestiae sed eveniet minus ullam quisquam."]