["Dolorum ducimus earum ullam omnis accusamus in in. Minus est non sequi sit est sunt voluptate. Adipisci aut ex et eveniet. Qui autem eveniet. Cupiditate illo exercitationem.", "Eum voluptatem deleniti iste accusantium assumenda nisi. Vel exercitationem deserunt consequuntur. Incidunt sed porro officia autem ut. Eos dicta vel voluptatem ab est necessitatibus. Necessitatibus sit quod consequatur facere vero aut iusto.", "Voluptates minima quidem fugit. Libero dolores optio et voluptatem. Facere maiores molestiae enim dolores. Perspiciatis nisi ullam tempore soluta ut. Velit ipsum unde ea voluptatem ipsam.", "Facere dicta rerum asperiores ipsam dolorum. Eum non voluptatem. Quidem harum recusandae.", "Qui velit modi. Aperiam rem temporibus debitis. Ea architecto velit quo fugit iusto. Ea fugiat vel unde recusandae possimus. Voluptatibus sunt quasi ad consequuntur omnis."]