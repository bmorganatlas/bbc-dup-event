["Perferendis tempore nam quis eum. Maxime reiciendis doloribus. Aliquid qui et accusamus dolor et. Repellat impedit ut corporis.", "Qui sit rerum numquam inventore placeat molestiae. Illo necessitatibus voluptatibus facilis dolorem expedita. Possimus mollitia ex expedita. Voluptatibus soluta enim molestiae quam.", "Perferendis aut quo. Nobis dolore consequatur. Est voluptas officia non cum qui. Assumenda deserunt optio qui fugit alias facere.", "Ad enim magnam. Asperiores sit deleniti est. Tempore id qui.", "Rerum qui quasi. Culpa nemo maiores laborum debitis qui qui voluptas. Qui voluptatem rem. Qui iste adipisci rerum aperiam sint debitis. Mollitia in autem consequatur alias quam atque est.", "Enim sint voluptas ea eius. Iure asperiores cupiditate. Distinctio asperiores ea autem porro in. Est facere beatae sed. Ducimus voluptas necessitatibus quia.", "Illo doloribus saepe ab. Non animi provident a. Enim sunt neque veritatis ad. Eligendi sint ab in sed quia placeat maiores. Aliquid rerum minima voluptatem qui voluptas.", "Est natus rerum. Animi et ut. Maxime autem recusandae ut soluta consectetur amet sit. Autem id dolor esse sit et.", "Quia quod cupiditate dolore est eum. Nulla incidunt fugit ducimus quae nesciunt quam. Est inventore pariatur exercitationem esse sed deserunt ipsum. Officia officiis sint nulla aliquid deleniti commodi.", "Accusantium iste ut consequatur est eum. Est veniam autem alias. Dolorem beatae accusantium dolores. Autem possimus culpa porro qui quia et aut."]