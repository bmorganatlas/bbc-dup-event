["Iure accusantium suscipit inventore rerum. Aut debitis id molestiae. Quas quis labore. Neque atque tempore rerum distinctio. Dolorem dolorum ut quam eligendi.", "Aut ea assumenda doloribus quidem nam praesentium facilis. Qui est distinctio. Quis beatae animi qui. Deleniti natus sapiente maxime quaerat sint ut nemo.", "Sunt est repellat praesentium atque quia inventore tempore. Est eos temporibus fugiat quis unde mollitia aut. Et culpa ut aut magni aliquid non odio. Voluptatem cumque qui iste sed omnis et esse.", "Unde illum omnis nam et deserunt. Dolorem voluptatem est ea quam explicabo necessitatibus. Quibusdam aut eum et nesciunt. Et vero ea minus.", "Quidem tempora nulla veritatis quaerat quo id enim. Vitae nobis dolor eos aut quis. Tempore sit non ut quod qui.", "Dolorem eum aut aliquam deleniti. Quisquam excepturi deserunt et. Praesentium aliquam id tenetur. Aut necessitatibus iure omnis ab.", "Consectetur qui autem veritatis. Qui optio nihil consequatur esse. Aliquam quia et blanditiis ex qui voluptatem est.", "Non in ratione corporis consectetur illum error. Eum facere sunt aliquid neque eveniet voluptatem ea. Est nobis placeat. Qui dolore hic sunt."]