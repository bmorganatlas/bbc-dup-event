["Occaecati quo aperiam voluptatem velit. Qui mollitia voluptatum. Quisquam sit maiores. Qui ex culpa voluptatem architecto.", "Ea et doloribus deserunt cum. Sint sit aperiam perspiciatis esse reprehenderit maiores ratione. Tempore maxime dicta nisi perferendis. Et quos incidunt ratione perferendis ipsam.", "Dolorem omnis minima facilis voluptas. Ratione et vitae aliquid nam asperiores nulla sit. Ullam omnis nesciunt sunt saepe et sint officiis. Odit voluptate iste consectetur.", "Tempora blanditiis debitis non sit. Labore in rerum ea doloribus. Dolores et sed qui eveniet qui repudiandae beatae. Voluptatum sed labore et. Minima rerum exercitationem.", "Occaecati sapiente ut hic debitis et iusto modi. Sed culpa libero consequuntur sunt voluptate cupiditate. Iusto tempore delectus corrupti. Aut voluptatibus maxime asperiores et dolorum. Quis nihil nam aperiam in.", "Iste sint qui dolorem dignissimos consequuntur. Aut laudantium sequi. Dolorem mollitia est distinctio non quia adipisci."]