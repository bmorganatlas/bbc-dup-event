["Quisquam quia maiores in modi. Tempore eos rerum id illo. Qui fuga vero ut. Aliquam dolor sit.", "Aperiam voluptates laboriosam eveniet ut itaque odit necessitatibus. Delectus ut voluptatem assumenda perferendis sit. Voluptas libero vero recusandae.", "Quam dolores distinctio doloribus voluptatem recusandae aut. Nemo ex debitis quae maiores dolores. Molestiae voluptatem voluptate sit nesciunt rerum. Soluta facilis quis fuga. Est qui ab."]