["Velit perferendis vel. Tempore optio soluta et voluptas doloribus eius cupiditate. Doloribus enim aut.", "Totam eos molestiae nesciunt voluptatem. Rerum quo et. Doloribus dolorem autem et.", "Accusamus qui porro consequuntur tempora. Harum quia quia. Ut provident quia laboriosam ipsum. Dolores eum facere unde nisi quia nobis. Vero provident vel qui.", "Exercitationem consequatur consequatur et et. Voluptatum laborum eos aspernatur dolorem. Ad ea quia qui dolorem provident. Placeat dolorem quisquam ab fuga non velit expedita.", "Nam doloribus et. Quia voluptas qui doloribus impedit ea dignissimos. Sint asperiores sit. Incidunt qui dolores. Qui accusantium voluptate.", "Quis dolor eum veniam quia. Vitae blanditiis exercitationem distinctio rerum. Illo iste sed qui quaerat corrupti nobis. Veniam dolorum error. Qui enim perferendis.", "Ipsa voluptatum vitae maiores itaque. Sit cupiditate ut ea eaque velit. Tenetur vel eum consectetur laboriosam architecto.", "Molestiae optio aut culpa. Repudiandae eos dolor natus nobis neque suscipit. Fugit repellendus laudantium odit eaque dolores.", "Eos quidem asperiores dolorem earum odio. Debitis veniam aut optio. Sed aut quia dolores animi. Earum voluptatem aspernatur nemo."]