["Voluptatem dolor tempore. Ratione adipisci itaque perferendis facere. Quia ut distinctio expedita dolor. Harum perferendis quis sit ex libero. Dolores illum quis non.", "Magni labore minus voluptas aliquam. Sint sequi aut illum. Ut non expedita repellat.", "Sed ab deserunt eligendi quaerat expedita dolorum dolores. Repudiandae reiciendis quo vitae molestiae nihil magnam est. Totam velit qui et. Est consequatur perspiciatis."]