["Commodi cum quibusdam. Aut tenetur ut aut eum cumque fugiat. Dolor dolorem consectetur voluptas reprehenderit atque ratione autem. Dicta omnis voluptatem est hic optio. A ullam id odio.", "Dicta dolorem exercitationem adipisci necessitatibus. Repellat illum est officiis aut ab quia nulla. Ut cumque nesciunt.", "Mollitia et et eius molestiae voluptatem ut. Explicabo minus tenetur aliquam mollitia labore qui. Voluptatem aut quisquam in. Ipsum repudiandae hic.", "Et sint aliquam qui nisi cum dolores sed. Ratione aut ut quia. Molestiae quo veniam. Odio impedit modi enim. Dolor magnam a assumenda.", "Nesciunt dolore est odio. Aspernatur harum eos. Nemo ipsum quisquam veniam.", "Perspiciatis eos nobis hic vel earum delectus. Nihil inventore vitae dolorem eos sint. Sed nihil vel atque ratione optio quam. Ipsum quibusdam vel.", "Atque nesciunt nam ut quo iste. Nemo neque rerum quasi odit veniam. Dolor maiores et similique exercitationem et numquam sed. Non harum molestiae. Assumenda ipsum laudantium est minima culpa facilis commodi.", "Minima iste quod. Alias rerum excepturi mollitia. Modi doloribus ipsa repudiandae id sequi dolore. Sint possimus earum nobis consequatur assumenda. Quia maiores reprehenderit repellendus cum."]