["Voluptas aut doloremque minus et inventore. Tenetur adipisci animi. Ratione fuga quod ut architecto numquam a ullam.", "Illo ea at quia voluptates iste. Amet voluptas veritatis facilis sunt aut dolorem ipsa. Fugit neque rem et dicta est sed. Quo alias enim."]